`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:46:19 11/04/2020
// Design Name: 
// Module Name:    test_VGA
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module test_VGA(
    input wire clk,           // board clock: 32 MHz quacho 100 MHz nexys4 
    input wire rst,         	// reset button

	// VGA input/output  
    output wire VGA_Hsync_n,  // horizontal sync output
    output wire VGA_Vsync_n,  // vertical sync output
    output wire [3:0] VGA_R,	// 4-bit VGA red output
    output wire [3:0] VGA_G,  // 4-bit VGA green output
    output wire [3:0] VGA_B,  // 4-bit VGA blue output
    output wire clkout,  
 	
	// input/output
	
	
	input wire bntr,
	input wire bntl
		
);

// TAMAÑO DE visualización 
parameter CAM_SCREEN_X = 184;
parameter CAM_SCREEN_Y = 184;

localparam AW = 6; // LOG2(CAM_SCREEN_X*CAM_SCREEN_Y)
localparam DW = 6;

// El color es RGB 222
localparam RED_VGA =   6'b110000;
localparam GREEN_VGA = 6'b001100;
localparam BLUE_VGA =  6'b000011;

// Clk 
wire clk12M;
wire clk25M;

// Conexión dual por ram

wire  [AW-1: 0] DP_RAM_addr_in;  
wire  [DW-1: 0] DP_RAM_data_in;
wire DP_RAM_regW;

reg  [AW-1: 0] DP_RAM_addr_out;  
	
// Conexión VGA Driver
wire [DW-1:0]data_mem;	   // Salida de dp_ram al driver VGA
wire [DW-1:0]data_RGB444;  // salida del driver VGA al puerto
wire [9:0]VGA_posX;		   // Determinar la pos de memoria que viene del VGA
wire [8:0]VGA_posY;		   // Determinar la pos de memoria que viene del VGA


/* ****************************************************************************
la pantalla VGA es RGB 444, pero el almacenamiento en memoria se hace 332
por lo tanto, los bits menos significactivos deben ser cero
**************************************************************************** */
	assign VGA_R = data_RGB444[5:4];
	assign VGA_G = data_RGB444[3:2];
	assign VGA_B = data_RGB444[1:0];



/* ****************************************************************************
  Este bloque se debe modificar según sea le caso. El ejemplo esta dado para
  fpga Spartan6 lx9 a 32MHz.
  usar "tools -> IP Generator ..."  y general el ip con Clocking Wizard
  el bloque genera un reloj de 25Mhz usado para el VGA , a partir de una frecuencia de 12 Mhz
**************************************************************************** */
assign clk12M =clk;

/*
cl_25_24_quartus clk25(
	.areset(rst),
	.inclk0(clk12M),
	.c0(clk25M)
	
);
*/
	reg [1:0] cfreq=0;
	assign clk25M = cfreq[0];
	always @(posedge clk) begin
			cfreq<=cfreq+1;
	end
assign clkout=clk25M;
/* ****************************************************************************
buffer_ram_dp buffer memoria dual port y reloj de lectura y escritura separados
Se debe configurar AW  según los calculos realizados en el Wp01
se recomiendia dejar DW a 8, con el fin de optimizar recursos  y hacer RGB 332
**************************************************************************** */
buffer_ram_dp #( AW,DW,"C:/Users/andre/Documents/GitHub/wp01-testvga-grupo-6/hdl/quartus/scr/image.men")
	DP_RAM(  
	.clk_w(clk25M), 
	.addr_in(DP_RAM_addr_in), 
	.data_in(DP_RAM_data_in),
	.regwrite(DP_RAM_regW), 
	.clk_r(clk25M), 
	.addr_out(DP_RAM_addr_out),
	.data_out(data_mem)
	);
	

/* ****************************************************************************
VGA_Driver640x480
**************************************************************************** */
VGA_Driver640x480 VGA640x480
(
	.rst(rst),
	.clk(clk25M), 				// 25MHz  para 60 hz de 640x480
	.pixelIn(data_mem), 		// entrada del valor de color  pixel RGB 444 
//	.pixelIn(RED_VGA), 		// entrada del valor de color  pixel RGB 444 
	.pixelOut(data_RGB444), // salida del valor pixel a la VGA 
	.Hsync_n(VGA_Hsync_n),	// señal de sincronizaciÓn en horizontal negada
	.Vsync_n(VGA_Vsync_n),	// señal de sincronizaciÓn en vertical negada 
	.posX(VGA_posX), 			// posición en horizontal del pixel siguiente
	.posY(VGA_posY) 			// posición en vertical  del pixel siguiente

);
 
/* ****************************************************************************
LÓgica para actualizar el pixel acorde con la buffer de memoria y el pixel de 
VGA si la imagen de la camara es menor que el display  VGA, los pixeles 
adicionales seran iguales al color del último pixel de memoria 
**************************************************************************** */

always @ (VGA_posX, VGA_posY) begin

		if ((VGA_posX<=160) && (VGA_posY<=120))
			DP_RAM_addr_out=0;
			
		else if ((VGA_posX<=320) && (VGA_posY<=120))
			DP_RAM_addr_out=16;
			
		else if ((VGA_posX<=480) && (VGA_posY<=120))
			DP_RAM_addr_out=55;
			
		else if ((VGA_posX<=640) && (VGA_posY<=120))
			DP_RAM_addr_out=40;
			
		else if ((VGA_posX<=160) && (VGA_posY<=240))
			DP_RAM_addr_out=1;
		
		else if ((VGA_posX<=320) && (VGA_posY<=240))
			DP_RAM_addr_out=12;
		
		else if ((VGA_posX<=480) && (VGA_posY<=240))
			DP_RAM_addr_out=52;
		
		else if ((VGA_posX<=640) && (VGA_posY<=240))
			DP_RAM_addr_out=17;
		
		else if ((VGA_posX<=160) && (VGA_posY<=360))
			DP_RAM_addr_out=34;
		
		else if ((VGA_posX<=320) && (VGA_posY<=360))
			DP_RAM_addr_out=46;
		
		else if ((VGA_posX<=480) && (VGA_posY<=360))
			DP_RAM_addr_out=5;
		
		else if ((VGA_posX<=640) && (VGA_posY<=360))
			DP_RAM_addr_out=30;
		
		else if ((VGA_posX<=160) && (VGA_posY<=480))
			DP_RAM_addr_out=0;
		
		else if ((VGA_posX<=320) && (VGA_posY<=480))
			DP_RAM_addr_out=15;
		
		else if ((VGA_posX<=480) && (VGA_posY<=480))
			DP_RAM_addr_out=24;
		
		else if ((VGA_posX<=640) && (VGA_posY<=480))
			DP_RAM_addr_out=63;

end

//assign DP_RAM_addr_out=10000;

/*****************************************************************************

este bloque debe crear un nuevo archivo 
**************************************************************************** */
 
 /*
 
 FSM_game  juego(
	 	.clk(clk25M),
		.rst(rst),
		.in1(btnr),
		.in2(btnr),
		.mem_px_addr(DP_RAM_addr_in),
		.mem_px_data(DP_RAM_data_in),
		.px_wr(DP_RAM_regW)
   );
	
	*/
endmodule
